`timescale 1ns / 1ps
//==============================================================================
// LeNet Layer 7 FC - Realistic RTL Test (Behavioral Model)
//
// Tests the first fully connected layer of LeNet-5:
//   Input:  (1, 256) - flattened from (1, 16, 4, 4)
//   Weight: (120, 256)
//   Output: (1, 120)
//
// GEMM: (1, 256) × (256, 120) → (1, 120)
//
// This testbench uses a behavioral model that performs the same
// tiled computation as the real RTL.
//
// Test vectors loaded from hex files generated by golden.py
//==============================================================================

module tb_lenet_layer7_fc;

    // Clock and timing
    parameter CLK_PERIOD = 10;
    parameter TIMEOUT_CYCLES = 50000;
    
    // GEMM dimensions
    parameter M = 1;        // Batch size
    parameter K = 256;      // Input features
    parameter N = 120;      // Output features
    parameter TILE = 8;     // Systolic array size
    
    // Derived tile counts
    parameter M_TILES = (M + TILE - 1) / TILE;  // 1
    parameter K_TILES = (K + TILE - 1) / TILE;  // 32
    parameter N_TILES = (N + TILE - 1) / TILE;  // 15
    
    reg clk = 0;
    always #(CLK_PERIOD/2) clk = ~clk;
    
    // =========================================================================
    // Test Data Storage
    // =========================================================================
    
    reg signed [7:0] A_mem [0:M*K-1];         // Input (1×256 = 256)
    reg signed [7:0] B_mem [0:K*N-1];         // Weights (256×120 = 30720)
    reg signed [31:0] C_expected [0:M*N-1];   // Expected output (1×120 = 120)
    reg signed [31:0] C_result [0:M*N-1];     // Result
    
    // =========================================================================
    // Behavioral Systolic Array Model
    // =========================================================================
    
    reg signed [31:0] pe_acc [0:TILE-1][0:TILE-1];
    reg signed [7:0] pe_weight [0:TILE-1][0:TILE-1];
    
    // =========================================================================
    // Test Variables
    // =========================================================================
    
    integer i, j, k;
    integer m_tile, n_tile, k_tile;
    integer m_start, n_start, k_start;
    integer m_size, k_size, n_size;
    integer cycle_count;
    integer tile_count;
    integer errors;
    integer total_compared;
    
    reg signed [7:0] a_val, b_val;
    reg signed [31:0] c_val, c_exp, diff;
    reg signed [31:0] mac_result;
    
    // =========================================================================
    // Helper Functions
    // =========================================================================
    
    function signed [7:0] get_A;
        input integer row, col;
    begin
        if (row < M && col < K)
            get_A = A_mem[row * K + col];
        else
            get_A = 8'sd0;
    end
    endfunction
    
    function signed [7:0] get_B;
        input integer row, col;
    begin
        if (row < K && col < N)
            get_B = B_mem[row * N + col];
        else
            get_B = 8'sd0;
    end
    endfunction
    
    // =========================================================================
    // Main Test
    // =========================================================================
    
    initial begin
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║      LeNet Layer 7 FC - Realistic RTL Test                       ║");
        $display("║      GEMM: (%0d, %0d) × (%0d, %0d) → (%0d, %0d)                          ║", M, K, K, N, M, N);
        $display("║      Tiled computation (%0d×%0d tiles)                               ║", TILE, TILE);
        $display("╚══════════════════════════════════════════════════════════════════╝");
        $display("");
        
        // Initialize
        cycle_count = 0;
        tile_count = 0;
        errors = 0;
        
        for (i = 0; i < M*N; i = i + 1) begin
            C_result[i] = 0;
        end
        
        // Load test vectors
        $display("[LOAD] Loading test vectors...");
        $readmemh("tests/realistic/lenet/test_vectors/layer7_input_int8.hex", A_mem);
        $readmemh("tests/realistic/lenet/test_vectors/layer7_weight_int8.hex", B_mem);
        $readmemh("tests/realistic/lenet/test_vectors/layer7_expected_int32.hex", C_expected);
        
        $display("  A[0]=%0d, A[1]=%0d", A_mem[0], A_mem[1]);
        $display("  B[0]=%0d, B[1]=%0d", B_mem[0], B_mem[1]);
        $display("  Expected C[0]=%0d, C[1]=%0d", C_expected[0], C_expected[1]);
        
        #(CLK_PERIOD*5);
        
        // Execute tiled GEMM
        $display("");
        $display("[EXEC] Starting tiled GEMM...");
        $display("  M=%0d, K=%0d, N=%0d", M, K, N);
        $display("  Tiles: M=%0d, K=%0d, N=%0d = %0d total", 
                 M_TILES, K_TILES, N_TILES, M_TILES * K_TILES * N_TILES);
        
        for (m_tile = 0; m_tile < M_TILES; m_tile = m_tile + 1) begin
            m_start = m_tile * TILE;
            m_size = ((m_start + TILE) > M) ? (M - m_start) : TILE;
            
            for (n_tile = 0; n_tile < N_TILES; n_tile = n_tile + 1) begin
                n_start = n_tile * TILE;
                n_size = ((n_start + TILE) > N) ? (N - n_start) : TILE;
                
                // Clear accumulators
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        pe_acc[i][j] = 0;
                    end
                end
                
                for (k_tile = 0; k_tile < K_TILES; k_tile = k_tile + 1) begin
                    k_start = k_tile * TILE;
                    k_size = ((k_start + TILE) > K) ? (K - k_start) : TILE;
                    
                    tile_count = tile_count + 1;
                    
                    // Load weights
                    for (i = 0; i < TILE; i = i + 1) begin
                        for (j = 0; j < TILE; j = j + 1) begin
                            pe_weight[i][j] = get_B(k_start + i, n_start + j);
                        end
                    end
                    cycle_count = cycle_count + TILE;
                    
                    // Compute MACs
                    for (k = 0; k < k_size; k = k + 1) begin
                        for (i = 0; i < m_size; i = i + 1) begin
                            a_val = get_A(m_start + i, k_start + k);
                            for (j = 0; j < n_size; j = j + 1) begin
                                b_val = pe_weight[k][j];
                                mac_result = $signed(a_val) * $signed(b_val);
                                pe_acc[i][j] = pe_acc[i][j] + mac_result;
                            end
                        end
                        cycle_count = cycle_count + 1;
                    end
                    
                    cycle_count = cycle_count + TILE;  // Drain
                    
                    if (tile_count % 100 == 0) begin
                        $display("  Tile %0d/%0d - %0d cycles",
                            tile_count, M_TILES * K_TILES * N_TILES, cycle_count);
                    end
                end
                
                // Write results
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        if (m_start + i < M && n_start + j < N) begin
                            C_result[(m_start + i) * N + (n_start + j)] = pe_acc[i][j];
                        end
                    end
                end
            end
        end
        
        $display("");
        $display("[DONE] GEMM complete: %0d tiles, %0d cycles", tile_count, cycle_count);
        
        // Verify
        $display("");
        $display("[VERIFY] Comparing results...");
        
        errors = 0;
        total_compared = 0;
        
        for (i = 0; i < M*N; i = i + 1) begin
            c_val = C_result[i];
            c_exp = C_expected[i];
            diff = (c_val > c_exp) ? (c_val - c_exp) : (c_exp - c_val);
            
            total_compared = total_compared + 1;
            
            if (diff > 0) begin
                errors = errors + 1;
                if (errors <= 10) begin
                    $display("  MISMATCH at [%0d]: got %0d, expected %0d", i, c_val, c_exp);
                end
            end
        end
        
        // Sample output
        $display("");
        $display("[SAMPLE] First 10 outputs:");
        for (i = 0; i < 10; i = i + 1) begin
            $display("  C[%0d] = %0d (expected %0d)", i, C_result[i], C_expected[i]);
        end
        
        // Summary
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║                      TEST SUMMARY                                ║");
        $display("╠══════════════════════════════════════════════════════════════════╣");
        $display("║  GEMM: (%0d × %0d) × (%0d × %0d) → (%0d × %0d)                            ║", M, K, K, N, M, N);
        $display("║  Tiles: %0d, Cycles: %0d                                       ║", tile_count, cycle_count);
        $display("║  Compared: %0d, Mismatches: %0d                                   ║", total_compared, errors);
        $display("╠══════════════════════════════════════════════════════════════════╣");
        
        if (errors == 0) begin
            $display("║  ✓ PASSED                                                       ║");
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER7 FC TEST PASSED! <<<");
        end else begin
            $display("║  ✗ FAILED: %0d mismatches                                       ║", errors);
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER7 FC TEST FAILED! <<<");
        end
        
        #(CLK_PERIOD * 10);
        $finish;
    end
    
    initial begin
        #(CLK_PERIOD * TIMEOUT_CYCLES);
        $display("ERROR: Timeout!");
        $finish;
    end

endmodule
