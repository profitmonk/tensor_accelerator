`timescale 1ns / 1ps
//==============================================================================
// Test: Multiple Sequential 4x4 GEMMs
// Validates system handles multiple back-to-back operations correctly
//==============================================================================
module tb_e2e_multi_gemm;
    parameter CLK = 10;
    parameter ARRAY_SIZE = 4;
    parameter SRAM_WIDTH = 256;

    reg clk = 0;
    reg rst_n = 0;
    always #(CLK/2) clk = ~clk;

    reg tpc_start = 0;
    reg [19:0] tpc_start_pc = 0;
    wire tpc_busy, tpc_done, tpc_error;
    reg global_sync_in = 0;
    wire sync_request;
    reg sync_grant = 0;
    reg [SRAM_WIDTH-1:0] noc_rx_data = 0;
    reg [19:0] noc_rx_addr = 0;
    reg noc_rx_valid = 0;
    wire noc_rx_ready;
    reg noc_rx_is_instr = 0;
    wire [SRAM_WIDTH-1:0] noc_tx_data;
    wire [19:0] noc_tx_addr;
    wire noc_tx_valid;
    reg noc_tx_ready = 1;
    wire [39:0] axi_awaddr, axi_araddr;
    wire [7:0] axi_awlen, axi_arlen;
    wire axi_awvalid, axi_arvalid, axi_wvalid, axi_wlast, axi_rready, axi_bready;
    wire [255:0] axi_wdata;
    reg axi_awready = 1, axi_arready = 1, axi_wready = 1;
    reg axi_bvalid = 0, axi_rvalid = 0, axi_rlast = 0;
    reg [1:0] axi_bresp = 0;
    reg [255:0] axi_rdata = 0;

    tensor_processing_cluster #(
        .ARRAY_SIZE(ARRAY_SIZE), .SRAM_WIDTH(SRAM_WIDTH),
        .SRAM_BANKS(4), .SRAM_DEPTH(256), .VPU_LANES(16)
    ) dut (
        .clk(clk), .rst_n(rst_n),
        .tpc_start(tpc_start), .tpc_start_pc(tpc_start_pc),
        .tpc_busy(tpc_busy), .tpc_done(tpc_done), .tpc_error(tpc_error),
        .global_sync_in(global_sync_in), .sync_request(sync_request), .sync_grant(sync_grant),
        .noc_rx_data(noc_rx_data), .noc_rx_addr(noc_rx_addr),
        .noc_rx_valid(noc_rx_valid), .noc_rx_ready(noc_rx_ready), .noc_rx_is_instr(noc_rx_is_instr),
        .noc_tx_data(noc_tx_data), .noc_tx_addr(noc_tx_addr),
        .noc_tx_valid(noc_tx_valid), .noc_tx_ready(noc_tx_ready),
        .axi_awaddr(axi_awaddr), .axi_awlen(axi_awlen), .axi_awvalid(axi_awvalid), .axi_awready(axi_awready),
        .axi_wdata(axi_wdata), .axi_wlast(axi_wlast), .axi_wvalid(axi_wvalid), .axi_wready(axi_wready),
        .axi_bresp(axi_bresp), .axi_bvalid(axi_bvalid), .axi_bready(axi_bready),
        .axi_araddr(axi_araddr), .axi_arlen(axi_arlen), .axi_arvalid(axi_arvalid), .axi_arready(axi_arready),
        .axi_rdata(axi_rdata), .axi_rlast(axi_rlast), .axi_rvalid(axi_rvalid), .axi_rready(axi_rready)
    );

    localparam OP_TENSOR = 8'h01;
    localparam OP_HALT = 8'hFF;

    // Two GEMMs: C1 = A1 × B1, C2 = A2 × B2
    // 
    // A1 = I (identity), B1 = [[1,2,3,4],[5,6,7,8],[9,10,11,12],[13,14,15,16]]
    // C1 = B1 (identity pass-through)
    //
    // A2 = [[2,0,0,0],[0,2,0,0],[0,0,2,0],[0,0,0,2]] (2×I)
    // B2 = [[1,1,1,1],[2,2,2,2],[3,3,3,3],[4,4,4,4]]
    // C2 = 2×B2 = [[2,2,2,2],[4,4,4,4],[6,6,6,6],[8,8,8,8]]

    reg [SRAM_WIDTH-1:0] row0, row1, row2, row3;
    integer i, errors;

    initial begin
        $display("");
        $display("╔════════════════════════════════════════════════════════════╗");
        $display("║         Multiple Sequential GEMM Test                      ║");
        $display("║         Two 4×4 GEMMs in one program                       ║");
        $display("╚════════════════════════════════════════════════════════════╝");
        
        //======================================================================
        // GEMM 1: C1 = I × B1 at addresses 0x00, 0x10, 0x20
        //======================================================================
        // B1^T (weights at 0x00)
        dut.sram_inst.bank_gen[0].bank_inst.mem[0] = {224'd0, 8'd13, 8'd9, 8'd5, 8'd1};
        dut.sram_inst.bank_gen[1].bank_inst.mem[0] = {224'd0, 8'd14, 8'd10, 8'd6, 8'd2};
        dut.sram_inst.bank_gen[2].bank_inst.mem[0] = {224'd0, 8'd15, 8'd11, 8'd7, 8'd3};
        dut.sram_inst.bank_gen[3].bank_inst.mem[0] = {224'd0, 8'd16, 8'd12, 8'd8, 8'd4};
        
        // A1 = I (activations at 0x10)
        dut.sram_inst.bank_gen[0].bank_inst.mem[4] = {224'd0, 8'd0, 8'd0, 8'd0, 8'd1};
        dut.sram_inst.bank_gen[1].bank_inst.mem[4] = {224'd0, 8'd0, 8'd0, 8'd1, 8'd0};
        dut.sram_inst.bank_gen[2].bank_inst.mem[4] = {224'd0, 8'd0, 8'd1, 8'd0, 8'd0};
        dut.sram_inst.bank_gen[3].bank_inst.mem[4] = {224'd0, 8'd1, 8'd0, 8'd0, 8'd0};

        //======================================================================
        // GEMM 2: C2 = 2I × B2 at addresses 0x40, 0x50, 0x60
        //======================================================================
        // B2^T (weights at 0x40 = word 16)
        dut.sram_inst.bank_gen[0].bank_inst.mem[16] = {224'd0, 8'd4, 8'd3, 8'd2, 8'd1};
        dut.sram_inst.bank_gen[1].bank_inst.mem[16] = {224'd0, 8'd4, 8'd3, 8'd2, 8'd1};
        dut.sram_inst.bank_gen[2].bank_inst.mem[16] = {224'd0, 8'd4, 8'd3, 8'd2, 8'd1};
        dut.sram_inst.bank_gen[3].bank_inst.mem[16] = {224'd0, 8'd4, 8'd3, 8'd2, 8'd1};
        
        // A2 = 2I (activations at 0x50 = word 20)
        dut.sram_inst.bank_gen[0].bank_inst.mem[20] = {224'd0, 8'd0, 8'd0, 8'd0, 8'd2};
        dut.sram_inst.bank_gen[1].bank_inst.mem[20] = {224'd0, 8'd0, 8'd0, 8'd2, 8'd0};
        dut.sram_inst.bank_gen[2].bank_inst.mem[20] = {224'd0, 8'd0, 8'd2, 8'd0, 8'd0};
        dut.sram_inst.bank_gen[3].bank_inst.mem[20] = {224'd0, 8'd2, 8'd0, 8'd0, 8'd0};

        //======================================================================
        // Program: GEMM1 → GEMM2 → HALT
        //======================================================================
        // GEMM1: dst=0x20, weights=0x00, acts=0x10
        dut.instr_mem[0] = {OP_TENSOR, 8'h01, 16'h0020, 16'h0010, 16'h0000, 16'd4, 16'd4, 16'd4, 16'd0};
        // GEMM2: dst=0x60, weights=0x40, acts=0x50
        dut.instr_mem[1] = {OP_TENSOR, 8'h01, 16'h0060, 16'h0050, 16'h0040, 16'd4, 16'd4, 16'd4, 16'd0};
        dut.instr_mem[2] = {OP_HALT, 120'd0};

        rst_n = 0; #(CLK*5); rst_n = 1; #(CLK*5);

        @(negedge clk); tpc_start = 1;
        @(posedge clk); @(posedge clk);
        @(negedge clk); tpc_start = 0;

        // Wait for completion (longer for 2 GEMMs)
        for (i = 0; i < 150; i = i + 1) begin
            @(posedge clk);
            if (tpc_done) i = 999;
        end
        #(CLK * 5);
        
        errors = 0;
        
        //======================================================================
        // Verify GEMM 1: C1 = B1 (output at 0x20 = word 8)
        //======================================================================
        $display("");
        $display("[GEMM 1] C1 = I × B1 (expect B1):");
        row0 = dut.sram_inst.bank_gen[0].bank_inst.mem[8];
        row1 = dut.sram_inst.bank_gen[1].bank_inst.mem[8];
        row2 = dut.sram_inst.bank_gen[2].bank_inst.mem[8];
        row3 = dut.sram_inst.bank_gen[3].bank_inst.mem[8];
        
        $display("  Row 0: [%0d,%0d,%0d,%0d] expect [1,2,3,4]",
            $signed(row0[31:0]), $signed(row0[63:32]), $signed(row0[95:64]), $signed(row0[127:96]));
        $display("  Row 1: [%0d,%0d,%0d,%0d] expect [5,6,7,8]",
            $signed(row1[31:0]), $signed(row1[63:32]), $signed(row1[95:64]), $signed(row1[127:96]));
        $display("  Row 2: [%0d,%0d,%0d,%0d] expect [9,10,11,12]",
            $signed(row2[31:0]), $signed(row2[63:32]), $signed(row2[95:64]), $signed(row2[127:96]));
        $display("  Row 3: [%0d,%0d,%0d,%0d] expect [13,14,15,16]",
            $signed(row3[31:0]), $signed(row3[63:32]), $signed(row3[95:64]), $signed(row3[127:96]));
        
        if (row0[31:0] != 1 || row0[63:32] != 2 || row0[95:64] != 3 || row0[127:96] != 4) errors = errors + 1;
        if (row1[31:0] != 5 || row1[63:32] != 6 || row1[95:64] != 7 || row1[127:96] != 8) errors = errors + 1;
        if (row2[31:0] != 9 || row2[63:32] != 10 || row2[95:64] != 11 || row2[127:96] != 12) errors = errors + 1;
        if (row3[31:0] != 13 || row3[63:32] != 14 || row3[95:64] != 15 || row3[127:96] != 16) errors = errors + 1;
        
        //======================================================================
        // Verify GEMM 2: C2 = 2×B2 (output at 0x60 = word 24)
        //======================================================================
        $display("");
        $display("[GEMM 2] C2 = 2I × B2 (expect 2×B2):");
        row0 = dut.sram_inst.bank_gen[0].bank_inst.mem[24];
        row1 = dut.sram_inst.bank_gen[1].bank_inst.mem[24];
        row2 = dut.sram_inst.bank_gen[2].bank_inst.mem[24];
        row3 = dut.sram_inst.bank_gen[3].bank_inst.mem[24];
        
        $display("  Row 0: [%0d,%0d,%0d,%0d] expect [2,2,2,2]",
            $signed(row0[31:0]), $signed(row0[63:32]), $signed(row0[95:64]), $signed(row0[127:96]));
        $display("  Row 1: [%0d,%0d,%0d,%0d] expect [4,4,4,4]",
            $signed(row1[31:0]), $signed(row1[63:32]), $signed(row1[95:64]), $signed(row1[127:96]));
        $display("  Row 2: [%0d,%0d,%0d,%0d] expect [6,6,6,6]",
            $signed(row2[31:0]), $signed(row2[63:32]), $signed(row2[95:64]), $signed(row2[127:96]));
        $display("  Row 3: [%0d,%0d,%0d,%0d] expect [8,8,8,8]",
            $signed(row3[31:0]), $signed(row3[63:32]), $signed(row3[95:64]), $signed(row3[127:96]));
        
        if (row0[31:0] != 2 || row0[63:32] != 2 || row0[95:64] != 2 || row0[127:96] != 2) errors = errors + 1;
        if (row1[31:0] != 4 || row1[63:32] != 4 || row1[95:64] != 4 || row1[127:96] != 4) errors = errors + 1;
        if (row2[31:0] != 6 || row2[63:32] != 6 || row2[95:64] != 6 || row2[127:96] != 6) errors = errors + 1;
        if (row3[31:0] != 8 || row3[63:32] != 8 || row3[95:64] != 8 || row3[127:96] != 8) errors = errors + 1;
        
        $display("");
        if (errors == 0) $display(">>> MULTI GEMM TEST PASSED! <<<");
        else $display(">>> MULTI GEMM TEST FAILED (%0d errors) <<<", errors);
        $finish;
    end
endmodule
