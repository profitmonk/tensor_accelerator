`timescale 1ns / 1ps
//==============================================================================
// LeNet Layer 3 Pool - Realistic RTL Test (Behavioral Model)
//
// Tests the first pooling layer of LeNet-5:
//   Input:  (1, 6, 24, 24) = 3456 elements
//   Output: (1, 6, 12, 12) = 864 elements
//   Operation: 2×2 average pooling
//
// Implementation:
//   For each 2×2 window: sum 4 values, shift right by 2 (divide by 4)
//
// Test vectors loaded from hex files generated by golden.py
//==============================================================================

module tb_lenet_layer3_pool;

    // Clock and timing
    parameter CLK_PERIOD = 10;
    parameter TIMEOUT_CYCLES = 50000;
    
    // Dimensions
    parameter IN_C = 6;
    parameter IN_H = 24;
    parameter IN_W = 24;
    parameter OUT_H = 12;
    parameter OUT_W = 12;
    parameter POOL_SIZE = 2;
    
    parameter IN_SIZE = IN_C * IN_H * IN_W;    // 3456
    parameter OUT_SIZE = IN_C * OUT_H * OUT_W; // 864
    
    reg clk = 0;
    always #(CLK_PERIOD/2) clk = ~clk;
    
    // =========================================================================
    // Test Data Storage
    // =========================================================================
    
    reg signed [7:0] input_mem [0:IN_SIZE-1];
    reg signed [7:0] expected_mem [0:OUT_SIZE-1];
    reg signed [7:0] result_mem [0:OUT_SIZE-1];
    
    // =========================================================================
    // Test Variables
    // =========================================================================
    
    integer c, oh, ow;
    integer in_idx, out_idx;
    integer cycle_count;
    integer errors;
    integer total_compared;
    
    reg signed [7:0] p00, p01, p10, p11;
    reg signed [15:0] sum;
    reg signed [7:0] avg;
    reg signed [7:0] expected_val, result_val;
    integer diff;
    
    // =========================================================================
    // Main Test
    // =========================================================================
    
    initial begin
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║      LeNet Layer 3 Pool - Realistic RTL Test                     ║");
        $display("║      Input: (%0d, %0d, %0d), Output: (%0d, %0d, %0d)                       ║", 
                 IN_C, IN_H, IN_W, IN_C, OUT_H, OUT_W);
        $display("║      2×2 Average Pooling                                         ║");
        $display("╚══════════════════════════════════════════════════════════════════╝");
        $display("");
        
        // Initialize
        cycle_count = 0;
        errors = 0;
        total_compared = 0;
        
        // Load test vectors
        $display("[LOAD] Loading test vectors...");
        $readmemh("tests/realistic/lenet/test_vectors/layer3_input_int8.hex", input_mem);
        $readmemh("tests/realistic/lenet/test_vectors/layer3_expected_int8.hex", expected_mem);
        
        $display("  Input[0]=%0d, Input[1]=%0d", input_mem[0], input_mem[1]);
        $display("  Expected[0]=%0d, Expected[1]=%0d", expected_mem[0], expected_mem[1]);
        
        #(CLK_PERIOD*5);
        
        // =====================================================================
        // Execute 2×2 Average Pooling
        // =====================================================================
        $display("");
        $display("[EXEC] Starting 2×2 average pooling...");
        $display("  Processing %0d channels × %0d×%0d output positions = %0d pools",
                 IN_C, OUT_H, OUT_W, OUT_SIZE);
        
        out_idx = 0;
        
        for (c = 0; c < IN_C; c = c + 1) begin
            for (oh = 0; oh < OUT_H; oh = oh + 1) begin
                for (ow = 0; ow < OUT_W; ow = ow + 1) begin
                    // Get 4 input values for this 2×2 window
                    // Input layout: [c, h, w] where c is slowest varying
                    p00 = input_mem[c * IN_H * IN_W + (oh*2 + 0) * IN_W + (ow*2 + 0)];
                    p01 = input_mem[c * IN_H * IN_W + (oh*2 + 0) * IN_W + (ow*2 + 1)];
                    p10 = input_mem[c * IN_H * IN_W + (oh*2 + 1) * IN_W + (ow*2 + 0)];
                    p11 = input_mem[c * IN_H * IN_W + (oh*2 + 1) * IN_W + (ow*2 + 1)];
                    
                    // Sum the 4 values
                    sum = $signed(p00) + $signed(p01) + $signed(p10) + $signed(p11);
                    
                    // Divide by 4 (arithmetic right shift by 2)
                    avg = sum >>> 2;
                    
                    // Store result
                    result_mem[out_idx] = avg;
                    out_idx = out_idx + 1;
                    
                    cycle_count = cycle_count + 1;
                end
            end
            
            // Progress per channel
            $display("  Channel %0d/%0d complete", c+1, IN_C);
        end
        
        $display("");
        $display("[DONE] Pooling complete: %0d output elements, %0d cycles", out_idx, cycle_count);
        
        // =====================================================================
        // Verify Results
        // =====================================================================
        $display("");
        $display("[VERIFY] Comparing results against expected...");
        
        errors = 0;
        total_compared = 0;
        
        for (out_idx = 0; out_idx < OUT_SIZE; out_idx = out_idx + 1) begin
            result_val = result_mem[out_idx];
            expected_val = expected_mem[out_idx];
            diff = (result_val > expected_val) ? (result_val - expected_val) : (expected_val - result_val);
            
            total_compared = total_compared + 1;
            
            // Allow ±1 tolerance for rounding differences
            if (diff > 1) begin
                errors = errors + 1;
                if (errors <= 10) begin
                    $display("  MISMATCH at [%0d]: got %0d, expected %0d (diff=%0d)",
                        out_idx, result_val, expected_val, diff);
                end
            end
        end
        
        // Print sample results
        $display("");
        $display("[SAMPLE] First 8 output values:");
        for (out_idx = 0; out_idx < 8; out_idx = out_idx + 1) begin
            $display("  Out[%0d] = %0d (expected %0d)", 
                     out_idx, result_mem[out_idx], expected_mem[out_idx]);
        end
        
        // =====================================================================
        // Summary
        // =====================================================================
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║                      TEST SUMMARY                                ║");
        $display("╠══════════════════════════════════════════════════════════════════╣");
        $display("║  Input:  (%0d, %0d, %0d) = %0d elements                              ║", IN_C, IN_H, IN_W, IN_SIZE);
        $display("║  Output: (%0d, %0d, %0d) = %0d elements                               ║", IN_C, OUT_H, OUT_W, OUT_SIZE);
        $display("║  Total cycles: %0d                                              ║", cycle_count);
        $display("║  Elements compared: %0d                                           ║", total_compared);
        $display("║  Mismatches (>1): %0d                                              ║", errors);
        $display("╠══════════════════════════════════════════════════════════════════╣");
        
        if (errors == 0) begin
            $display("║  ✓ PASSED: All outputs within tolerance                        ║");
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER3 POOL TEST PASSED! <<<");
        end else begin
            $display("║  ✗ FAILED: %0d mismatches found                                 ║", errors);
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER3 POOL TEST FAILED! <<<");
        end
        
        $display("");
        #(CLK_PERIOD * 10);
        $finish;
    end
    
    // Timeout
    initial begin
        #(CLK_PERIOD * TIMEOUT_CYCLES);
        $display("ERROR: Timeout!");
        $finish;
    end

endmodule
