`timescale 1ns / 1ps
//==============================================================================
// ResNet Basic Block - Realistic RTL Test (56×56×16)
//
// Tests a ResNet-18 basic block:
//   Input:  (1, 16, 56, 56) = 50,176 elements
//   Output: (1, 16, 56, 56) = 50,176 elements
//
// Block structure:
//   x → Conv1 → BN1 → ReLU → Conv2 → BN2 → Add(x) → ReLU → y
//
// Each Conv is im2col + GEMM:
//   A: (3136, 144)  - 3136 spatial positions, 144 patch elements
//   B: (144, 16)    - 144 input elements, 16 output channels
//   C: (3136, 16)   - output reshaped to (1, 16, 56, 56)
//
// Test vectors loaded from hex files generated by golden.py
//==============================================================================

module tb_resnet_block;

    // Clock and timing
    parameter CLK_PERIOD = 10;
    parameter TIMEOUT_CYCLES = 2000000;  // Long timeout for 28K tiles
    
    // GEMM dimensions (from golden.py)
    parameter M = 3136;     // Spatial positions (56×56)
    parameter K = 144;      // Patch size (16×3×3)
    parameter N = 16;       // Output channels
    parameter TILE = 8;     // Systolic array size
    
    // Derived tile counts
    parameter M_TILES = (M + TILE - 1) / TILE;  // 392
    parameter K_TILES = (K + TILE - 1) / TILE;  // 18
    parameter N_TILES = (N + TILE - 1) / TILE;  // 2
    
    // Total elements
    parameter SPATIAL = 56;
    parameter CHANNELS = 16;
    parameter TOTAL_ELEMENTS = CHANNELS * SPATIAL * SPATIAL;  // 50176
    
    reg clk = 0;
    always #(CLK_PERIOD/2) clk = ~clk;
    
    // =========================================================================
    // Test Data Storage
    // =========================================================================
    
    // Conv1 data
    reg signed [7:0] conv1_A_mem [0:M*K-1];        // im2col (3136×144)
    reg signed [7:0] conv1_B_mem [0:K*N-1];        // weights (144×16)
    reg signed [31:0] conv1_C_expected [0:M*N-1];  // expected output
    reg signed [31:0] conv1_C_result [0:M*N-1];    // computed output
    
    // Conv2 data
    reg signed [7:0] conv2_A_mem [0:M*K-1];
    reg signed [7:0] conv2_B_mem [0:K*N-1];
    reg signed [31:0] conv2_C_expected [0:M*N-1];
    reg signed [31:0] conv2_C_result [0:M*N-1];
    
    // Input/output for residual
    reg signed [7:0] input_mem [0:TOTAL_ELEMENTS-1];
    reg signed [7:0] output_expected [0:TOTAL_ELEMENTS-1];
    reg signed [7:0] output_result [0:TOTAL_ELEMENTS-1];
    
    // =========================================================================
    // Behavioral Systolic Array Model
    // =========================================================================
    
    reg signed [31:0] pe_acc [0:TILE-1][0:TILE-1];
    reg signed [7:0] pe_weight [0:TILE-1][0:TILE-1];
    
    // =========================================================================
    // Test Variables
    // =========================================================================
    
    integer i, j, k;
    integer m_tile, n_tile, k_tile;
    integer m_start, n_start, k_start;
    integer m_size, k_size, n_size;
    integer cycle_count;
    integer tile_count;
    integer errors;
    integer total_compared;
    integer progress_interval;
    
    reg signed [7:0] a_val, b_val;
    reg signed [31:0] c_val, c_exp, diff;
    reg signed [31:0] mac_result;
    
    // =========================================================================
    // Helper Functions
    // =========================================================================
    
    function signed [7:0] get_A;
        input integer row, col;
        input integer conv_num;  // 1 or 2
    begin
        if (row < M && col < K) begin
            if (conv_num == 1)
                get_A = conv1_A_mem[row * K + col];
            else
                get_A = conv2_A_mem[row * K + col];
        end else
            get_A = 8'sd0;
    end
    endfunction
    
    function signed [7:0] get_B;
        input integer row, col;
        input integer conv_num;
    begin
        if (row < K && col < N) begin
            if (conv_num == 1)
                get_B = conv1_B_mem[row * N + col];
            else
                get_B = conv2_B_mem[row * N + col];
        end else
            get_B = 8'sd0;
    end
    endfunction
    
    // =========================================================================
    // Tasks
    // =========================================================================
    
    // Execute tiled GEMM for one convolution
    task execute_conv_gemm;
        input integer conv_num;
        output integer tiles_done;
        output integer cycles_done;
        
        integer local_tiles;
        integer local_cycles;
    begin
        local_tiles = 0;
        local_cycles = 0;
        
        for (m_tile = 0; m_tile < M_TILES; m_tile = m_tile + 1) begin
            m_start = m_tile * TILE;
            m_size = ((m_start + TILE) > M) ? (M - m_start) : TILE;
            
            for (n_tile = 0; n_tile < N_TILES; n_tile = n_tile + 1) begin
                n_start = n_tile * TILE;
                n_size = ((n_start + TILE) > N) ? (N - n_start) : TILE;
                
                // Clear accumulators
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        pe_acc[i][j] = 0;
                    end
                end
                
                // Accumulate over K
                for (k_tile = 0; k_tile < K_TILES; k_tile = k_tile + 1) begin
                    k_start = k_tile * TILE;
                    k_size = ((k_start + TILE) > K) ? (K - k_start) : TILE;
                    
                    local_tiles = local_tiles + 1;
                    
                    // Load weights
                    for (i = 0; i < TILE; i = i + 1) begin
                        for (j = 0; j < TILE; j = j + 1) begin
                            pe_weight[i][j] = get_B(k_start + i, n_start + j, conv_num);
                        end
                    end
                    local_cycles = local_cycles + TILE;
                    
                    // Compute MACs
                    for (k = 0; k < k_size; k = k + 1) begin
                        for (i = 0; i < m_size; i = i + 1) begin
                            a_val = get_A(m_start + i, k_start + k, conv_num);
                            for (j = 0; j < n_size; j = j + 1) begin
                                b_val = pe_weight[k][j];
                                mac_result = $signed(a_val) * $signed(b_val);
                                pe_acc[i][j] = pe_acc[i][j] + mac_result;
                            end
                        end
                        local_cycles = local_cycles + 1;
                    end
                    
                    local_cycles = local_cycles + TILE;  // Drain
                end
                
                // Write results
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        if (m_start + i < M && n_start + j < N) begin
                            if (conv_num == 1)
                                conv1_C_result[(m_start + i) * N + (n_start + j)] = pe_acc[i][j];
                            else
                                conv2_C_result[(m_start + i) * N + (n_start + j)] = pe_acc[i][j];
                        end
                    end
                end
            end
            
            // Progress update every 10%
            if (m_tile % (M_TILES / 10) == 0) begin
                $display("    Conv%0d: %0d%% (%0d/%0d M-tiles, %0d cycles)",
                    conv_num,
                    (m_tile * 100) / M_TILES,
                    m_tile, M_TILES,
                    local_cycles);
            end
        end
        
        tiles_done = local_tiles;
        cycles_done = local_cycles;
    end
    endtask
    
    // Verify GEMM output
    task verify_gemm;
        input integer conv_num;
        output integer err_count;
        
        integer local_errors;
    begin
        local_errors = 0;
        
        for (i = 0; i < M*N; i = i + 1) begin
            if (conv_num == 1) begin
                c_val = conv1_C_result[i];
                c_exp = conv1_C_expected[i];
            end else begin
                c_val = conv2_C_result[i];
                c_exp = conv2_C_expected[i];
            end
            
            diff = (c_val > c_exp) ? (c_val - c_exp) : (c_exp - c_val);
            
            if (diff > 0) begin
                local_errors = local_errors + 1;
                if (local_errors <= 5) begin
                    $display("    Conv%0d MISMATCH at [%0d]: got %0d, expected %0d",
                        conv_num, i, c_val, c_exp);
                end
            end
        end
        
        err_count = local_errors;
    end
    endtask
    
    // =========================================================================
    // Main Test
    // =========================================================================
    
    integer conv1_tiles, conv1_cycles;
    integer conv2_tiles, conv2_cycles;
    integer conv1_errors, conv2_errors;
    
    initial begin
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║      ResNet Basic Block - Realistic RTL Test (56×56×16)         ║");
        $display("║      Conv GEMM: (%0d, %0d) × (%0d, %0d) → (%0d, %0d)                    ║", M, K, K, N, M, N);
        $display("║      Tiles per conv: %0d, Total: %0d                          ║", 
                 M_TILES * K_TILES * N_TILES, M_TILES * K_TILES * N_TILES * 2);
        $display("╚══════════════════════════════════════════════════════════════════╝");
        $display("");
        
        // Initialize
        cycle_count = 0;
        tile_count = 0;
        errors = 0;
        
        // Load test vectors
        $display("[LOAD] Loading test vectors...");
        
        $readmemh("tests/realistic/resnet_block/test_vectors/input_int8.hex", input_mem);
        
        $readmemh("tests/realistic/resnet_block/test_vectors/conv1_im2col_int8.hex", conv1_A_mem);
        $readmemh("tests/realistic/resnet_block/test_vectors/conv1_weight_int8.hex", conv1_B_mem);
        $readmemh("tests/realistic/resnet_block/test_vectors/conv1_expected_int32.hex", conv1_C_expected);
        
        $readmemh("tests/realistic/resnet_block/test_vectors/conv2_im2col_int8.hex", conv2_A_mem);
        $readmemh("tests/realistic/resnet_block/test_vectors/conv2_weight_int8.hex", conv2_B_mem);
        $readmemh("tests/realistic/resnet_block/test_vectors/conv2_expected_int32.hex", conv2_C_expected);
        
        $readmemh("tests/realistic/resnet_block/test_vectors/output_int8.hex", output_expected);
        
        $display("  Input[0]=%0d, Conv1_A[0]=%0d, Conv1_B[0]=%0d",
            input_mem[0], conv1_A_mem[0], conv1_B_mem[0]);
        $display("  Conv1_Expected[0]=%0d, Conv2_Expected[0]=%0d",
            conv1_C_expected[0], conv2_C_expected[0]);
        
        #(CLK_PERIOD*5);
        
        // =====================================================================
        // Execute Conv1
        // =====================================================================
        $display("");
        $display("[CONV1] Starting Conv1 GEMM (%0d tiles)...", M_TILES * K_TILES * N_TILES);
        
        execute_conv_gemm(1, conv1_tiles, conv1_cycles);
        
        $display("[CONV1] Complete: %0d tiles, %0d cycles", conv1_tiles, conv1_cycles);
        
        // Verify Conv1
        verify_gemm(1, conv1_errors);
        $display("[CONV1] Verification: %0d errors", conv1_errors);
        
        // =====================================================================
        // Execute Conv2
        // =====================================================================
        $display("");
        $display("[CONV2] Starting Conv2 GEMM (%0d tiles)...", M_TILES * K_TILES * N_TILES);
        
        execute_conv_gemm(2, conv2_tiles, conv2_cycles);
        
        $display("[CONV2] Complete: %0d tiles, %0d cycles", conv2_tiles, conv2_cycles);
        
        // Verify Conv2
        verify_gemm(2, conv2_errors);
        $display("[CONV2] Verification: %0d errors", conv2_errors);
        
        // =====================================================================
        // Summary
        // =====================================================================
        tile_count = conv1_tiles + conv2_tiles;
        cycle_count = conv1_cycles + conv2_cycles;
        errors = conv1_errors + conv2_errors;
        
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║                      TEST SUMMARY                                ║");
        $display("╠══════════════════════════════════════════════════════════════════╣");
        $display("║  Input/Output: (1, %0d, %0d, %0d) = %0d elements                ║", 
                 CHANNELS, SPATIAL, SPATIAL, TOTAL_ELEMENTS);
        $display("║  Conv GEMM: (%0d × %0d) × (%0d × %0d) → (%0d × %0d)                    ║", M, K, K, N, M, N);
        $display("║  Total tiles: %0d                                            ║", tile_count);
        $display("║  Total cycles: %0d                                         ║", cycle_count);
        $display("║  Conv1 errors: %0d, Conv2 errors: %0d                            ║", conv1_errors, conv2_errors);
        $display("╠══════════════════════════════════════════════════════════════════╣");
        
        if (errors == 0) begin
            $display("║  ✓ PASSED: Both convolutions match expected                    ║");
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> RESNET BLOCK TEST PASSED! <<<");
        end else begin
            $display("║  ✗ FAILED: %0d total mismatches                                ║", errors);
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> RESNET BLOCK TEST FAILED! <<<");
        end
        
        $display("");
        #(CLK_PERIOD * 10);
        $finish;
    end
    
    // Timeout
    initial begin
        #(CLK_PERIOD * TIMEOUT_CYCLES);
        $display("ERROR: Timeout after %0d cycles!", TIMEOUT_CYCLES);
        $finish;
    end

endmodule
