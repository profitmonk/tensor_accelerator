`timescale 1ns / 1ps
//==============================================================================
// LeNet Layer 1 Conv - Realistic RTL Test (Behavioral Model)
//
// Tests the first convolution layer of LeNet-5:
//   Input:  (1, 1, 28, 28) 
//   Weight: (6, 1, 5, 5)
//   Output: (1, 6, 24, 24)
//
// Computation via im2col + GEMM:
//   A: (576, 25)  - im2col transformed input patches
//   B: (25, 6)    - reshaped weights
//   C: (576, 6)   - output (reshape to 24×24×6)
//
// This testbench uses a behavioral systolic array model that performs
// the same tiled computation as the real RTL, verifying the dataflow
// and comparing against Python golden model outputs.
//
// Test vectors loaded from hex files generated by golden.py
//==============================================================================

module tb_lenet_layer1_conv;

    // Clock and timing
    parameter CLK_PERIOD = 10;
    parameter TIMEOUT_CYCLES = 100000;
    
    // GEMM dimensions (from golden.py)
    parameter M = 576;      // Number of patches (24×24)
    parameter K = 25;       // Patch size (1×5×5)
    parameter N = 6;        // Output channels
    parameter TILE = 8;     // Systolic array size
    
    // Derived tile counts
    parameter M_TILES = (M + TILE - 1) / TILE;  // 72
    parameter K_TILES = (K + TILE - 1) / TILE;  // 4 (with padding)
    parameter N_TILES = (N + TILE - 1) / TILE;  // 1 (with padding)
    
    reg clk = 0;
    always #(CLK_PERIOD/2) clk = ~clk;
    
    // =========================================================================
    // Test Data Storage
    // =========================================================================
    
    // Input matrices (loaded from hex files)
    reg signed [7:0] A_mem [0:M*K-1];         // im2col input (576×25 = 14400)
    reg signed [7:0] B_mem [0:K*N-1];         // weights (25×6 = 150)
    reg signed [31:0] C_expected [0:M*N-1];   // expected output (576×6 = 3456)
    
    // Output accumulator
    reg signed [31:0] C_result [0:M*N-1];
    
    // =========================================================================
    // Behavioral Systolic Array Model
    // Performs 8×8 tiled GEMM identical to RTL
    // =========================================================================
    
    // PE accumulators (8×8 grid)
    reg signed [31:0] pe_acc [0:TILE-1][0:TILE-1];
    reg signed [7:0] pe_weight [0:TILE-1][0:TILE-1];
    
    // =========================================================================
    // Test Variables
    // =========================================================================
    
    integer i, j, k, t;
    integer m_tile, n_tile, k_tile;
    integer m_start, m_end, n_start, n_end, k_start, k_end;
    integer m_size, k_size, n_size;
    integer cycle_count;
    integer tile_count;
    integer errors;
    integer total_compared;
    
    reg signed [7:0] a_val, b_val;
    reg signed [31:0] c_val, c_exp;
    reg signed [31:0] diff;
    reg signed [31:0] mac_result;
    
    // =========================================================================
    // Helper Functions
    // =========================================================================
    
    // Get A matrix element with bounds checking
    function signed [7:0] get_A;
        input integer row, col;
    begin
        if (row < M && col < K)
            get_A = A_mem[row * K + col];
        else
            get_A = 8'sd0;
    end
    endfunction
    
    // Get B matrix element with bounds checking  
    function signed [7:0] get_B;
        input integer row, col;
    begin
        if (row < K && col < N)
            get_B = B_mem[row * N + col];
        else
            get_B = 8'sd0;
    end
    endfunction
    
    // =========================================================================
    // Main Test
    // =========================================================================
    
    initial begin
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║      LeNet Layer 1 Conv - Realistic RTL Test                     ║");
        $display("║      GEMM: (%0d, %0d) × (%0d, %0d) → (%0d, %0d)                            ║", M, K, K, N, M, N);
        $display("║      Tiled computation (%0d×%0d tiles)                               ║", TILE, TILE);
        $display("╚══════════════════════════════════════════════════════════════════╝");
        $display("");
        
        // Initialize
        cycle_count = 0;
        tile_count = 0;
        errors = 0;
        total_compared = 0;
        
        // Initialize output accumulator
        for (i = 0; i < M*N; i = i + 1) begin
            C_result[i] = 0;
        end
        
        // Load test vectors
        $display("[LOAD] Loading test vectors from hex files...");
        $readmemh("tests/realistic/lenet/test_vectors/layer1_im2col_int8.hex", A_mem);
        $readmemh("tests/realistic/lenet/test_vectors/layer1_weight_int8.hex", B_mem);
        $readmemh("tests/realistic/lenet/test_vectors/layer1_expected_int32.hex", C_expected);
        
        // Verify load
        $display("  A[0]=%0d, A[1]=%0d, A[2]=%0d", A_mem[0], A_mem[1], A_mem[2]);
        $display("  B[0]=%0d, B[1]=%0d, B[2]=%0d", B_mem[0], B_mem[1], B_mem[2]);
        $display("  Expected C[0]=%0d, C[1]=%0d", C_expected[0], C_expected[1]);
        
        #(CLK_PERIOD*5);
        
        // =====================================================================
        // Execute Tiled GEMM (Output-Stationary)
        // For each output tile (m, n), accumulate across all k tiles
        // =====================================================================
        $display("");
        $display("[EXEC] Starting tiled GEMM...");
        $display("  M=%0d, K=%0d, N=%0d", M, K, N);
        $display("  Tiles: M=%0d, K=%0d, N=%0d", M_TILES, K_TILES, N_TILES);
        $display("  Total tile operations: %0d", M_TILES * K_TILES * N_TILES);
        $display("");
        
        for (m_tile = 0; m_tile < M_TILES; m_tile = m_tile + 1) begin
            m_start = m_tile * TILE;
            m_size = ((m_start + TILE) > M) ? (M - m_start) : TILE;
            
            for (n_tile = 0; n_tile < N_TILES; n_tile = n_tile + 1) begin
                n_start = n_tile * TILE;
                n_size = ((n_start + TILE) > N) ? (N - n_start) : TILE;
                
                // Clear PE accumulators for this output tile
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        pe_acc[i][j] = 0;
                    end
                end
                
                // Accumulate across K dimension
                for (k_tile = 0; k_tile < K_TILES; k_tile = k_tile + 1) begin
                    k_start = k_tile * TILE;
                    k_size = ((k_start + TILE) > K) ? (K - k_start) : TILE;
                    
                    tile_count = tile_count + 1;
                    
                    // Load weights into PE array
                    for (i = 0; i < TILE; i = i + 1) begin
                        for (j = 0; j < TILE; j = j + 1) begin
                            pe_weight[i][j] = get_B(k_start + i, n_start + j);
                        end
                    end
                    cycle_count = cycle_count + TILE;  // Weight load cycles
                    
                    // Compute: each PE does MAC for its position
                    // This models the systolic dataflow
                    for (k = 0; k < k_size; k = k + 1) begin
                        for (i = 0; i < m_size; i = i + 1) begin
                            a_val = get_A(m_start + i, k_start + k);
                            for (j = 0; j < n_size; j = j + 1) begin
                                b_val = pe_weight[k][j];
                                mac_result = $signed(a_val) * $signed(b_val);
                                pe_acc[i][j] = pe_acc[i][j] + mac_result;
                            end
                        end
                        cycle_count = cycle_count + 1;
                    end
                    
                    // Drain cycles
                    cycle_count = cycle_count + TILE;
                end
                
                // Write accumulated results to output
                for (i = 0; i < TILE; i = i + 1) begin
                    for (j = 0; j < TILE; j = j + 1) begin
                        if (m_start + i < M && n_start + j < N) begin
                            C_result[(m_start + i) * N + (n_start + j)] = pe_acc[i][j];
                        end
                    end
                end
                
                // Progress update every 10 M-tiles
                if (m_tile % 10 == 0 && n_tile == 0 && tile_count > 0) begin
                    $display("  Progress: M-tile %0d/%0d, %0d tiles done, %0d cycles",
                        m_tile, M_TILES, tile_count, cycle_count);
                end
            end
        end
        
        $display("");
        $display("[DONE] GEMM complete: %0d tiles, %0d cycles", tile_count, cycle_count);
        
        // =====================================================================
        // Verify Results
        // =====================================================================
        $display("");
        $display("[VERIFY] Comparing results against expected...");
        
        errors = 0;
        total_compared = 0;
        
        for (i = 0; i < M; i = i + 1) begin
            for (j = 0; j < N; j = j + 1) begin
                c_val = C_result[i * N + j];
                c_exp = C_expected[i * N + j];
                diff = (c_val > c_exp) ? (c_val - c_exp) : (c_exp - c_val);
                
                total_compared = total_compared + 1;
                
                if (diff > 0) begin
                    errors = errors + 1;
                    if (errors <= 10) begin
                        $display("  MISMATCH at [%0d,%0d]: got %0d, expected %0d (diff=%0d)",
                            i, j, c_val, c_exp, diff);
                    end
                end
            end
        end
        
        // Print sample results
        $display("");
        $display("[SAMPLE] First 5 output values:");
        for (i = 0; i < 5; i = i + 1) begin
            $display("  C[%0d] = %0d (expected %0d)", i, C_result[i], C_expected[i]);
        end
        
        $display("");
        $display("[SAMPLE] Last 5 output values:");
        for (i = M*N-5; i < M*N; i = i + 1) begin
            $display("  C[%0d] = %0d (expected %0d)", i, C_result[i], C_expected[i]);
        end
        
        // =====================================================================
        // Summary
        // =====================================================================
        $display("");
        $display("╔══════════════════════════════════════════════════════════════════╗");
        $display("║                      TEST SUMMARY                                ║");
        $display("╠══════════════════════════════════════════════════════════════════╣");
        $display("║  GEMM: (%0d × %0d) × (%0d × %0d) → (%0d × %0d)                            ║", M, K, K, N, M, N);
        $display("║  Tiles executed: %0d                                            ║", tile_count);
        $display("║  Total cycles: %0d                                           ║", cycle_count);
        $display("║  Elements compared: %0d                                        ║", total_compared);
        $display("║  Mismatches: %0d                                                 ║", errors);
        $display("╠══════════════════════════════════════════════════════════════════╣");
        
        if (errors == 0) begin
            $display("║  ✓ PASSED: All outputs match expected values                   ║");
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER1 CONV TEST PASSED! <<<");
        end else begin
            $display("║  ✗ FAILED: %0d mismatches found                                 ║", errors);
            $display("╚══════════════════════════════════════════════════════════════════╝");
            $display("");
            $display(">>> LENET LAYER1 CONV TEST FAILED! <<<");
        end
        
        $display("");
        #(CLK_PERIOD * 10);
        $finish;
    end
    
    // Timeout watchdog
    initial begin
        #(CLK_PERIOD * TIMEOUT_CYCLES);
        $display("");
        $display("ERROR: Test timeout after %0d cycles!", TIMEOUT_CYCLES);
        $display(">>> LENET LAYER1 CONV TEST FAILED (TIMEOUT)! <<<");
        $finish;
    end

endmodule
